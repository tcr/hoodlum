module Main (
);
endmodule

